netcdf LMDZ_stdpressurelevels {
dimensions:
	LMDZ_STDPRESSURELEVELS = 17 ;
	LMDZ_STDPRESSURELEVELSedges = 18 ;
variables:
	double LMDZ_STDPRESSURELEVELS(LMDZ_STDPRESSURELEVELS) ;
		LMDZ_STDPRESSURELEVELS:units = "mb" ;
		LMDZ_STDPRESSURELEVELS:positive = "down" ;
		LMDZ_STDPRESSURELEVELS:point_spacing = "uneven" ;
		LMDZ_STDPRESSURELEVELS:edges = "LMDZ_STDPRESSURELEVELSedges" ;
	double LMDZ_STDPRESSURELEVELSedges(LMDZ_STDPRESSURELEVELSedges) ;
		LMDZ_STDPRESSURELEVELSedges:edges = " " ;
data:

 LMDZ_STDPRESSURELEVELS = 10, 20, 30, 50, 70, 100, 150, 200, 250, 300, 400, 
    500, 600, 700, 850, 925, 1000 ;

 LMDZ_STDPRESSURELEVELSedges = 5, 15, 25, 40, 60, 85, 125, 175, 225, 275, 
    350, 450, 550, 650, 775, 887.5, 962.5, 1037.5 ;
}
