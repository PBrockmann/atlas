netcdf ECMWF50_stdpressurelevels {
dimensions:
	ECMWF50_STDPRESSURELEVELS = 50 ;
	ECMWF50_STDPRESSURELEVELSedges = 51 ;
variables:
	double ECMWF50_STDPRESSURELEVELS(ECMWF50_STDPRESSURELEVELS) ;
		ECMWF50_STDPRESSURELEVELS:units = "mb" ;
		ECMWF50_STDPRESSURELEVELS:positive = "down" ;
		ECMWF50_STDPRESSURELEVELS:point_spacing = "uneven" ;
		ECMWF50_STDPRESSURELEVELS:edges = "ECMWF50_STDPRESSURELEVELSedges" ;
	double ECMWF50_STDPRESSURELEVELSedges(ECMWF50_STDPRESSURELEVELSedges) ;
		ECMWF50_STDPRESSURELEVELSedges:edges = " " ;
data:

 ECMWF50_STDPRESSURELEVELS = 
0.100000, 0.316500, 0.593200, 0.952100, 1.384900, 1.889000, 2.469500, 3.140700, 3.928500, 4.876100, 6.041300, 7.485100, 9.273800, 11.490100, 14.235900, 17.638000, 21.853000, 27.075400, 33.545800, 41.562400, 51.494900, 63.487500, 77.579800, 93.837200, 112.267400, 132.940400, 155.898300, 181.154400, 208.649400, 238.325800, 270.153000, 304.046500, 339.889100, 377.546600, 416.878900, 457.744200, 500.000000, 543.496900, 588.068400, 633.514400, 679.579800, 725.928500, 772.110200, 817.524200, 861.375600, 902.628700, 939.952000, 971.660900, 995.653300, 1009.339600 ;

 ECMWF50_STDPRESSURELEVELSedges = 
0.000000, 0.200100, 0.433000, 0.753500, 1.150800, 1.619000, 2.159000, 2.780100, 3.501400, 4.355600, 5.396500, 6.686200, 8.284000, 10.263700, 12.716400, 15.755400, 19.520500, 24.185500, 29.965300, 37.126300, 45.998600, 56.991100, 69.983900, 85.175800, 102.498700, 122.036200, 143.844600, 167.951900, 194.356800, 222.942000, 253.709600, 286.596400, 321.496600, 358.281500, 396.811800, 436.945900, 478.542500, 521.457500, 565.536400, 610.600500, 656.428300, 702.731500, 749.125500, 795.094900, 839.953400, 882.798000, 922.459400, 957.444700, 985.877300, 1005.429200, 1013.250000 ;

}
